// 4 Bit Full Adder

module FourBitFullAdder(A, B, C, carry, sum);
    input [3:0] A, [3:0] B, C;
    output carry, sum;
    reg carry, sum;

